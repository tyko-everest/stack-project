`ifndef _consts_h
`define _consts_h

localparam DATA_STACK_SIZE = 8;
localparam RET_STACK_SIZE = 8;
localparam STACK_WIDTH = 8;
localparam PROG_MEM_SIZE = 16;
localparam PROG_MEM_WIDTH = 4;

`endif
